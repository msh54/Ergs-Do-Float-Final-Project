module counter(start_count1,start_count2,end_count,start_recovery, start_ref1, start_ref2, end_ref3, end_recovery,clk,reset);
input  clk,start_drive,start_recovery, start_ref1, start_ref2, end_ref3, end_recovery;
output[31:0] start_count1,start_count2,end_count;


endmodule
