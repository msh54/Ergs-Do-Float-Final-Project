module processor_testbench;

endmodule