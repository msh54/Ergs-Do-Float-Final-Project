module rusher(rush,start_recovery, start_ref1, start_ref2, end_ref3, end_recovery,clk);


endmodule
