
module ratioer(ratio,start_drive,start_recovery,count_clock);
	input start_drive, start_recovery,count_clock;
	output[31:0] ratio;
	wire[31:0] recovery_count,drive_count,divResult;


	wire reset;
	counter _counter(drive_count,recovery_count,start_drive,start_recovery,count_clock);
	// counter(drive_count,recovery_count,start_drive,start_recovery,clk);
	
	//wire divResult;
	
	divider _div(recovery_count,drive_count,divResult);
	
	
	// In counter, there is a 5 cycle delay between enable and reset; can use ratio != 0, because the numerator 0 will be reset to 0
	assign enable = start_drive && (reset != 0) && (divResult != 0);
	
	register _ratReg(.clk(count_clock), .in_en(enable), .data_in(divResult), .data_out(ratio), .clr(1'b0));

endmodule

/*
Have a counter adding at a certain rate, either incrementing drive or recovery

every time start_drive is high, on the positive edge, calculate the ratio


*/ 