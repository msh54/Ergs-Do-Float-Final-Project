module exor(out,in1,in2);
	input in1,in2;
	output out;
	xor _xor(out,in1,in2);
endmodule
